// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus II Version 15.0.0 Build 145 04/22/2015 SJ Web Edition
// Created on Thu Oct 27 17:09:32 2016

// synthesis message_off 10175

`timescale 1ns/1ns

module SM1 (
    reset,clock,x0,x1);

    input reset;
    input clock;
    input x0;
    input x1;
    tri0 reset;
    tri0 x0;
    tri0 x1;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter state1=0,state2=1,state3=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or x0 or x1)
    begin
        if (reset) begin
            reg_fstate <= state1;
        end
        else begin
            case (fstate)
                state1: begin
                    if ((x0 & ~(x1)))
                        reg_fstate <= state2;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;
                end
                state2: begin
                    if (~(x1))
                        reg_fstate <= state1;
                    else if (x1)
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;
                end
                state3: begin
                    if ((~(x1) & ~(x0)))
                        reg_fstate <= state1;
                    else if ((x1 | x0))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;
                end
                default: begin
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // SM1
