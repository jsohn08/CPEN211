module cpu(reset, clk);


endmodule;
