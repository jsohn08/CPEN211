module cpu_tb();
  reg 
